** Generated for: hspiceD
** Generated on: Dec  1 03:58:12 2023
** Design library name: cad4
** Design cell name: lfsr
** Design view name: schematic
.GLOBAL vdd! vss!


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_bip
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_dio
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_dio_33
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_mim
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_dio_dnw
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_dio_18
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_bip_npn
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_33
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_rfrtmom
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_mos_cap_25
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_18
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_disres
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_res
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_dio_na
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_rfmos_33
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_dio_hvt
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_rfmvar
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_rfmos_18
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_na
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_dio_na33
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_dio_lvt
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_rfres_sa
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_na33
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_dio_esd
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_rfmim
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_dio_25od33
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_25od33
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_mos_cap
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_dio_25
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_dio_25ud18
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_25
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_rfmos
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_25ud18
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_dio_na25od33
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_rfjvar
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_rfmos_25
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_rtmom
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_na25od33
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_dio_na25
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_rfres_rpo
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_hvt
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_rfind
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_rfmvar_25
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_na25
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65RF/1.0c/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt_lvt

** Library name: cad2
** Cell name: INVD1
** View name: schematic
.subckt INVD1 vi vo
m0 vo vi vdd! vdd! pch l=60e-9 w=400e-9 m=1 nf=1 sd=200e-9 ad=70e-15 as=70e-15 pd=1.15e-6 ps=1.15e-6 nrd=250e-3 nrs=250e-3 sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m1 vo vi vss! vss! nch l=60e-9 w=300e-9 m=1 nf=1 sd=200e-9 ad=52.5e-15 as=52.5e-15 pd=950e-9 ps=950e-9 nrd=333.333e-3 nrs=333.333e-3 sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
.ends INVD1
** End of subcircuit definition.

** Library name: cad3
** Cell name: NAND2_balanced
** View name: schematic
.subckt NAND2_balanced a b out
mpmos1 out b vdd! vdd! pch l=60e-9 w=450e-9 m=1 nf=1 sd=200e-9 ad=78.75e-15 as=78.75e-15 pd=1.25e-6 ps=1.25e-6 nrd=222.222e-3 nrs=222.222e-3 sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
mpmos0 out a vdd! vdd! pch l=60e-9 w=450e-9 m=1 nf=1 sd=200e-9 ad=78.75e-15 as=78.75e-15 pd=1.25e-6 ps=1.25e-6 nrd=222.222e-3 nrs=222.222e-3 sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
mnmos1 net14 b vss! vss! nch l=60e-9 w=350e-9 m=1 nf=1 sd=200e-9 ad=61.25e-15 as=61.25e-15 pd=1.05e-6 ps=1.05e-6 nrd=285.714e-3 nrs=285.714e-3 sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
mnmos0 out a net14 vss! nch l=60e-9 w=350e-9 m=1 nf=1 sd=200e-9 ad=61.25e-15 as=61.25e-15 pd=1.05e-6 ps=1.05e-6 nrd=285.714e-3 nrs=285.714e-3 sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
.ends NAND2_balanced
** End of subcircuit definition.

** Library name: cad4
** Cell name: NOR
** View name: schematic
.subckt NOR a b z
m1 z a net15 vdd! pch l=60e-9 w=450e-9 m=1 nf=1 sd=200e-9 ad=78.75e-15 as=78.75e-15 pd=1.25e-6 ps=1.25e-6 nrd=222.222e-3 nrs=222.222e-3 sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m0 net15 b vdd! vdd! pch l=60e-9 w=450e-9 m=1 nf=1 sd=200e-9 ad=78.75e-15 as=78.75e-15 pd=1.25e-6 ps=1.25e-6 nrd=222.222e-3 nrs=222.222e-3 sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m3 z b vss! vss! nch l=60e-9 w=350e-9 m=1 nf=1 sd=200e-9 ad=61.25e-15 as=61.25e-15 pd=1.05e-6 ps=1.05e-6 nrd=285.714e-3 nrs=285.714e-3 sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m2 z a vss! vss! nch l=60e-9 w=350e-9 m=1 nf=1 sd=200e-9 ad=61.25e-15 as=61.25e-15 pd=1.05e-6 ps=1.05e-6 nrd=285.714e-3 nrs=285.714e-3 sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
.ends NOR
** End of subcircuit definition.

** Library name: cad4
** Cell name: CLK
** View name: schematic
.subckt CLK clk clki clki_bar
xi1 clki_bar clki INVD1
xi0 clk clki_bar INVD1
.ends CLK
** End of subcircuit definition.

** Library name: cad4
** Cell name: RST
** View name: schematic
.subckt RST rst rst_bar
xi0 rst rst_bar INVD1
.ends RST
** End of subcircuit definition.

** Library name: cad4
** Cell name: GATE
** View name: schematic
.subckt GATE a a_bar vi vo
m0 vi a vo vdd! pch l=60e-9 w=350e-9 m=1 nf=1 sd=200e-9 ad=61.25e-15 as=61.25e-15 pd=1.05e-6 ps=1.05e-6 nrd=285.714e-3 nrs=285.714e-3 sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m1 vi a_bar vo vss! nch l=60e-9 w=300e-9 m=1 nf=1 sd=200e-9 ad=52.5e-15 as=52.5e-15 pd=950e-9 ps=950e-9 nrd=333.333e-3 nrs=333.333e-3 sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
.ends GATE
** End of subcircuit definition.

** Library name: cad4
** Cell name: DFSR
** View name: schematic
.subckt DFSR clk d q rst
xi3 net016 net033 INVD1
xi13 net033 q INVD1
xi1 net9 net13 INVD1
xi0 d net7 INVD1
xi12 net024 net13 net17 NAND2_balanced
xi6 net033 rst net019 NOR
xi8 clk net020 net028 CLK
xi9 rst net024 RST
xi17 net028 net020 net9 net17 GATE
xi16 net028 net020 net13 net016 GATE
xi15 net020 net028 net016 net019 GATE
xi14 net020 net028 net7 net9 GATE
.ends DFSR
** End of subcircuit definition.

** Library name: cad4
** Cell name: XOR2
** View name: schematic
.subckt XOR2 a b z
xi3 net20 net19 z NAND2_balanced
xi2 net11 b net19 NAND2_balanced
xi1 a net11 net20 NAND2_balanced
xi0 a b net11 NAND2_balanced
.ends XOR2
** End of subcircuit definition.

** Library name: cad4
** Cell name: XOR4
** View name: schematic
.subckt XOR4 a b c d z
xi12 a b net7 XOR2
xi13 c d net6 XOR2
xi14 net7 net6 z XOR2
.ends XOR4
** End of subcircuit definition.

** Library name: cad4
** Cell name: OR
** View name: schematic
.subckt OR a b z
xi0 net7 z INVD1
xi1 a b net7 NOR
.ends OR
** End of subcircuit definition.

** Library name: cad4
** Cell name: lfsr
** View name: schematic
xi15 clk state<1> state<0> rst DFSR
xi14 clk state<2> state<1> rst DFSR
xi13 clk state<3> state<2> rst DFSR
xi12 clk state<4> state<3> rst DFSR
xi11 clk state<5> state<4> rst DFSR
xi10 clk state<6> state<5> rst DFSR
xi9 clk state<7> state<6> rst DFSR
xi8 clk state<8> state<7> rst DFSR
xi7 clk state<9> state<8> rst DFSR
xi6 clk state<10> state<9> rst DFSR
xi5 clk state<11> state<10> rst DFSR
xi4 clk state<12> state<11> rst DFSR
xi3 clk state<13> state<12> rst DFSR
xi2 clk state<14> state<13> rst DFSR
xi1 clk state<15> state<14> rst DFSR
xi0 clk net064 state<15> vss! DFSR
xi23 state<0> state<2> state<3> state<5> net069 XOR4
xi22 net069 rst net064 OR
.END
